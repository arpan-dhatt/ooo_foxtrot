// Logical functional unit

module fu_logical (
    fu_if.fu fu
);

  // Empty module body

endmodule
